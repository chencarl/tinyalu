class tinyalu_config extends uvm_object;
    `uvm_object_utils(tinyalu_config)
    
    function new(string name = "");
        super.new(name);
    endfunction
endclass